----------------------------------------------------------------------------------
-- Design Name   : led_top
-- Create Date   : 2015/12/31
-- Module Name   : 
-- Project Name  : 
-- Target Devices: 
-- Tool Versions : 
-- Description   : 
-- Revision      :
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
--The MIT License (MIT)
--
--Copyright (c) 2015 
--
--Permission is hereby granted, free of charge, to any person obtaining a copy
--of this software and associated documentation files (the "Software"), to deal
--in the Software without restriction, including without limitation the rights
--to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--copies of the Software, and to permit persons to whom the Software is
--furnished to do so, subject to the following conditions:
--
--The above copyright notice and this permission notice shall be included in all
--copies or substantial portions of the Software.
--
--THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--SOFTWARE.
----------------------------------------------------------------------------------



-- Library Define
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;





entity niosii_top is
    Port ( 
		p_clk_50Mhz		: in  std_logic;    	
		
		p_button		: in  std_logic_vector( 1 downto 0 );
		p_led_out		: out std_logic_vector( 7 downto 0 );
		
		p_pwm_dir       : out std_logic_vector(1 downto 0);
		p_pwm_out       : out std_logic_vector(1 downto 0);
		
		p_uart_0_rxd    : in  std_logic;
		p_uart_0_txd    : out std_logic;				
		
		p_epcs_flash_dclk	 : out std_logic;                           
		p_epcs_flash_sce	 : out std_logic;                           
		p_epcs_flash_sdo	 : out std_logic;                          
		p_epcs_flash_data0 	 : in  std_logic
		
		);
end niosii_top;


architecture Behavioral of niosii_top is


    component niosii is
        port (
            clk_clk                          : in  std_logic                    := 'X'; -- clk
            pio_0_external_connection_export : out std_logic_vector(7 downto 0);        -- export
            reset_reset_n                    : in  std_logic                    := 'X'; -- reset_n
            uart_0_rxd                       : in  std_logic                    := 'X'; -- rxd
            uart_0_txd                       : out std_logic;                           -- txd
            ip_pwm_dir                       : out std_logic_vector(1 downto 0);        -- dir
            ip_pwm_out                       : out std_logic_vector(1 downto 0);        -- out			
            epcs_flash_dclk                  : out std_logic;                           -- dclk
            epcs_flash_sce                   : out std_logic;                           -- sce
            epcs_flash_sdo                   : out std_logic;                           -- sdo
            epcs_flash_data0                 : in  std_logic                    := 'X'  -- data0			
        );
    end component niosii;


		
	signal s_reset_n			: std_logic;
begin

	s_reset_n <= p_button(0);
	

    u0 : component niosii
        port map (
            clk_clk                          => p_clk_50Mhz,
            pio_0_external_connection_export => p_led_out,
            reset_reset_n                    => s_reset_n,
            uart_0_rxd                       => p_uart_0_rxd, 
            uart_0_txd                       => p_uart_0_txd,  
            ip_pwm_dir                       => p_pwm_dir,
            ip_pwm_out                       => p_pwm_out,			
            epcs_flash_dclk                  => p_epcs_flash_dclk,
            epcs_flash_sce                   => p_epcs_flash_sce,
            epcs_flash_sdo                   => p_epcs_flash_sdo,
            epcs_flash_data0                 => p_epcs_flash_data0			
        );	
		
end Behavioral;
