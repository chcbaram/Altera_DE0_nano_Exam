-- altera_epcq_controller_core.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity altera_epcq_controller_core is
	generic (
		DEVICE_FAMILY     : string  := "Cyclone IV E";
		ADDR_WIDTH        : integer := 19;
		ASMI_ADDR_WIDTH   : integer := 24;
		ASI_WIDTH         : integer := 1;
		CS_WIDTH          : integer := 1;
		CHIP_SELS         : integer := 1;
		ENABLE_4BYTE_ADDR : integer := 0
	);
	port (
		clk                  : in  std_logic                     := '0';             --          clock_sink.clk
		reset_n              : in  std_logic                     := '0';             --               reset.reset_n
		avl_csr_read         : in  std_logic                     := '0';             --             avl_csr.read
		avl_csr_waitrequest  : out std_logic;                                        --                    .waitrequest
		avl_csr_write        : in  std_logic                     := '0';             --                    .write
		avl_csr_addr         : in  std_logic_vector(2 downto 0)  := (others => '0'); --                    .address
		avl_csr_wrdata       : in  std_logic_vector(31 downto 0) := (others => '0'); --                    .writedata
		avl_csr_rddata       : out std_logic_vector(31 downto 0);                    --                    .readdata
		avl_csr_rddata_valid : out std_logic;                                        --                    .readdatavalid
		avl_mem_write        : in  std_logic                     := '0';             --             avl_mem.write
		avl_mem_burstcount   : in  std_logic_vector(6 downto 0)  := (others => '0'); --                    .burstcount
		avl_mem_waitrequest  : out std_logic;                                        --                    .waitrequest
		avl_mem_read         : in  std_logic                     := '0';             --                    .read
		avl_mem_addr         : in  std_logic_vector(18 downto 0) := (others => '0'); --                    .address
		avl_mem_wrdata       : in  std_logic_vector(31 downto 0) := (others => '0'); --                    .writedata
		avl_mem_rddata       : out std_logic_vector(31 downto 0);                    --                    .readdata
		avl_mem_rddata_valid : out std_logic;                                        --                    .readdatavalid
		avl_mem_byteenable   : in  std_logic_vector(3 downto 0)  := (others => '0'); --                    .byteenable
		asmi_status_out      : in  std_logic_vector(7 downto 0)  := (others => '0'); --     asmi_status_out.conduit_status_out
		asmi_epcs_id         : in  std_logic_vector(7 downto 0)  := (others => '0'); --        asmi_epcs_id.conduit_epcs_id
		asmi_illegal_erase   : in  std_logic                     := '0';             --  asmi_illegal_erase.conduit_illegal_erase
		asmi_illegal_write   : in  std_logic                     := '0';             --  asmi_illegal_write.conduit_illegal_write
		ddasi_dataoe         : in  std_logic_vector(0 downto 0)  := (others => '0'); --        ddasi_dataoe.conduit_ddasi_dataoe
		ddasi_dclk           : in  std_logic                     := '0';             --          ddasi_dclk.conduit_ddasi_dclk
		ddasi_scein          : in  std_logic_vector(0 downto 0)  := (others => '0'); --         ddasi_scein.conduit_ddasi_scein
		ddasi_sdoin          : in  std_logic_vector(0 downto 0)  := (others => '0'); --         ddasi_sdoin.conduit_ddasi_sdoin
		asmi_busy            : in  std_logic                     := '0';             --           asmi_busy.conduit_busy
		asmi_data_valid      : in  std_logic                     := '0';             --     asmi_data_valid.conduit_data_valid
		asmi_dataout         : in  std_logic_vector(7 downto 0)  := (others => '0'); --        asmi_dataout.conduit_dataout
		epcq_dataout         : in  std_logic_vector(0 downto 0)  := (others => '0'); --        epcq_dataout.conduit_epcq_dataout
		ddasi_dataout        : out std_logic_vector(0 downto 0);                     --       ddasi_dataout.conduit_ddasi_dataout
		asmi_read_rdid       : out std_logic;                                        --      asmi_read_rdid.conduit_read_rdid
		asmi_read_status     : out std_logic;                                        --    asmi_read_status.conduit_read_status
		asmi_read_sid        : out std_logic;                                        --       asmi_read_sid.conduit_read_sid
		asmi_bulk_erase      : out std_logic;                                        --     asmi_bulk_erase.conduit_bulk_erase
		asmi_sector_erase    : out std_logic;                                        --   asmi_sector_erase.conduit_sector_erase
		asmi_sector_protect  : out std_logic;                                        -- asmi_sector_protect.conduit_sector_protect
		epcq_dclk            : out std_logic;                                        --           epcq_dclk.conduit_epcq_dclk
		epcq_scein           : out std_logic_vector(0 downto 0);                     --          epcq_scein.conduit_epcq_scein
		epcq_sdoin           : out std_logic_vector(0 downto 0);                     --          epcq_sdoin.conduit_epcq_sdoin
		epcq_dataoe          : out std_logic_vector(0 downto 0);                     --         epcq_dataoe.conduit_epcq_dataoe
		asmi_clkin           : out std_logic;                                        --          asmi_clkin.conduit_clkin
		asmi_reset           : out std_logic;                                        --          asmi_reset.conduit_reset
		asmi_sce             : out std_logic_vector(0 downto 0);                     --            asmi_sce.conduit_asmi_sce
		asmi_addr            : out std_logic_vector(23 downto 0);                    --           asmi_addr.conduit_addr
		asmi_datain          : out std_logic_vector(7 downto 0);                     --         asmi_datain.conduit_datain
		asmi_fast_read       : out std_logic;                                        --      asmi_fast_read.conduit_fast_read
		asmi_rden            : out std_logic;                                        --           asmi_rden.conduit_rden
		asmi_shift_bytes     : out std_logic;                                        --    asmi_shift_bytes.conduit_shift_bytes
		asmi_wren            : out std_logic;                                        --           asmi_wren.conduit_wren
		asmi_write           : out std_logic;                                        --          asmi_write.conduit_write
		asmi_rdid_out        : in  std_logic_vector(7 downto 0)  := (others => '0'); --       asmi_rdid_out.conduit_rdid_out
		asmi_en4b_addr       : out std_logic;                                        --      asmi_en4b_addr.conduit_en4b_addr
		irq                  : out std_logic                                         --    interrupt_sender.irq
	);
end entity altera_epcq_controller_core;

architecture rtl of altera_epcq_controller_core is
	component altera_epcq_controller_arb is
		generic (
			DEVICE_FAMILY     : string  := "";
			ADDR_WIDTH        : integer := 19;
			ASMI_ADDR_WIDTH   : integer := 24;
			ASI_WIDTH         : integer := 1;
			CS_WIDTH          : integer := 1;
			CHIP_SELS         : integer := 1;
			ENABLE_4BYTE_ADDR : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset_n              : in  std_logic                     := 'X';             -- reset_n
			avl_csr_read         : in  std_logic                     := 'X';             -- read
			avl_csr_waitrequest  : out std_logic;                                        -- waitrequest
			avl_csr_write        : in  std_logic                     := 'X';             -- write
			avl_csr_addr         : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avl_csr_wrdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_csr_rddata       : out std_logic_vector(31 downto 0);                    -- readdata
			avl_csr_rddata_valid : out std_logic;                                        -- readdatavalid
			avl_mem_write        : in  std_logic                     := 'X';             -- write
			avl_mem_burstcount   : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			avl_mem_waitrequest  : out std_logic;                                        -- waitrequest
			avl_mem_read         : in  std_logic                     := 'X';             -- read
			avl_mem_addr         : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			avl_mem_wrdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_mem_rddata       : out std_logic_vector(31 downto 0);                    -- readdata
			avl_mem_rddata_valid : out std_logic;                                        -- readdatavalid
			avl_mem_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			asmi_status_out      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- conduit_status_out
			asmi_epcs_id         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- conduit_epcs_id
			asmi_illegal_erase   : in  std_logic                     := 'X';             -- conduit_illegal_erase
			asmi_illegal_write   : in  std_logic                     := 'X';             -- conduit_illegal_write
			ddasi_dataoe         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- conduit_ddasi_dataoe
			ddasi_dclk           : in  std_logic                     := 'X';             -- conduit_ddasi_dclk
			ddasi_scein          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- conduit_ddasi_scein
			ddasi_sdoin          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- conduit_ddasi_sdoin
			asmi_busy            : in  std_logic                     := 'X';             -- conduit_busy
			asmi_data_valid      : in  std_logic                     := 'X';             -- conduit_data_valid
			asmi_dataout         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- conduit_dataout
			epcq_dataout         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- conduit_epcq_dataout
			ddasi_dataout        : out std_logic_vector(0 downto 0);                     -- conduit_ddasi_dataout
			asmi_read_rdid       : out std_logic;                                        -- conduit_read_rdid
			asmi_read_status     : out std_logic;                                        -- conduit_read_status
			asmi_read_sid        : out std_logic;                                        -- conduit_read_sid
			asmi_bulk_erase      : out std_logic;                                        -- conduit_bulk_erase
			asmi_sector_erase    : out std_logic;                                        -- conduit_sector_erase
			asmi_sector_protect  : out std_logic;                                        -- conduit_sector_protect
			epcq_dclk            : out std_logic;                                        -- conduit_epcq_dclk
			epcq_scein           : out std_logic_vector(0 downto 0);                     -- conduit_epcq_scein
			epcq_sdoin           : out std_logic_vector(0 downto 0);                     -- conduit_epcq_sdoin
			epcq_dataoe          : out std_logic_vector(0 downto 0);                     -- conduit_epcq_dataoe
			asmi_clkin           : out std_logic;                                        -- conduit_clkin
			asmi_reset           : out std_logic;                                        -- conduit_reset
			asmi_sce             : out std_logic_vector(0 downto 0);                     -- conduit_asmi_sce
			asmi_addr            : out std_logic_vector(23 downto 0);                    -- conduit_addr
			asmi_datain          : out std_logic_vector(7 downto 0);                     -- conduit_datain
			asmi_fast_read       : out std_logic;                                        -- conduit_fast_read
			asmi_rden            : out std_logic;                                        -- conduit_rden
			asmi_shift_bytes     : out std_logic;                                        -- conduit_shift_bytes
			asmi_wren            : out std_logic;                                        -- conduit_wren
			asmi_write           : out std_logic;                                        -- conduit_write
			asmi_rdid_out        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- conduit_rdid_out
			asmi_en4b_addr       : out std_logic;                                        -- conduit_en4b_addr
			irq                  : out std_logic                                         -- irq
		);
	end component altera_epcq_controller_arb;

begin

	device_family_check : if DEVICE_FAMILY /= "Cyclone IV E" generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	addr_width_check : if ADDR_WIDTH /= 19 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	asmi_addr_width_check : if ASMI_ADDR_WIDTH /= 24 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	asi_width_check : if ASI_WIDTH /= 1 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	cs_width_check : if CS_WIDTH /= 1 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	chip_sels_check : if CHIP_SELS /= 1 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	enable_4byte_addr_check : if ENABLE_4BYTE_ADDR /= 0 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	altera_epcq_controller_core : component altera_epcq_controller_arb
		generic map (
			DEVICE_FAMILY     => "Cyclone IV E",
			ADDR_WIDTH        => 19,
			ASMI_ADDR_WIDTH   => 24,
			ASI_WIDTH         => 1,
			CS_WIDTH          => 1,
			CHIP_SELS         => 1,
			ENABLE_4BYTE_ADDR => 0
		)
		port map (
			clk                  => clk,                  --          clock_sink.clk
			reset_n              => reset_n,              --               reset.reset_n
			avl_csr_read         => avl_csr_read,         --             avl_csr.read
			avl_csr_waitrequest  => avl_csr_waitrequest,  --                    .waitrequest
			avl_csr_write        => avl_csr_write,        --                    .write
			avl_csr_addr         => avl_csr_addr,         --                    .address
			avl_csr_wrdata       => avl_csr_wrdata,       --                    .writedata
			avl_csr_rddata       => avl_csr_rddata,       --                    .readdata
			avl_csr_rddata_valid => avl_csr_rddata_valid, --                    .readdatavalid
			avl_mem_write        => avl_mem_write,        --             avl_mem.write
			avl_mem_burstcount   => avl_mem_burstcount,   --                    .burstcount
			avl_mem_waitrequest  => avl_mem_waitrequest,  --                    .waitrequest
			avl_mem_read         => avl_mem_read,         --                    .read
			avl_mem_addr         => avl_mem_addr,         --                    .address
			avl_mem_wrdata       => avl_mem_wrdata,       --                    .writedata
			avl_mem_rddata       => avl_mem_rddata,       --                    .readdata
			avl_mem_rddata_valid => avl_mem_rddata_valid, --                    .readdatavalid
			avl_mem_byteenable   => avl_mem_byteenable,   --                    .byteenable
			asmi_status_out      => asmi_status_out,      --     asmi_status_out.conduit_status_out
			asmi_epcs_id         => asmi_epcs_id,         --        asmi_epcs_id.conduit_epcs_id
			asmi_illegal_erase   => asmi_illegal_erase,   --  asmi_illegal_erase.conduit_illegal_erase
			asmi_illegal_write   => asmi_illegal_write,   --  asmi_illegal_write.conduit_illegal_write
			ddasi_dataoe         => ddasi_dataoe,         --        ddasi_dataoe.conduit_ddasi_dataoe
			ddasi_dclk           => ddasi_dclk,           --          ddasi_dclk.conduit_ddasi_dclk
			ddasi_scein          => ddasi_scein,          --         ddasi_scein.conduit_ddasi_scein
			ddasi_sdoin          => ddasi_sdoin,          --         ddasi_sdoin.conduit_ddasi_sdoin
			asmi_busy            => asmi_busy,            --           asmi_busy.conduit_busy
			asmi_data_valid      => asmi_data_valid,      --     asmi_data_valid.conduit_data_valid
			asmi_dataout         => asmi_dataout,         --        asmi_dataout.conduit_dataout
			epcq_dataout         => epcq_dataout,         --        epcq_dataout.conduit_epcq_dataout
			ddasi_dataout        => ddasi_dataout,        --       ddasi_dataout.conduit_ddasi_dataout
			asmi_read_rdid       => asmi_read_rdid,       --      asmi_read_rdid.conduit_read_rdid
			asmi_read_status     => asmi_read_status,     --    asmi_read_status.conduit_read_status
			asmi_read_sid        => asmi_read_sid,        --       asmi_read_sid.conduit_read_sid
			asmi_bulk_erase      => asmi_bulk_erase,      --     asmi_bulk_erase.conduit_bulk_erase
			asmi_sector_erase    => asmi_sector_erase,    --   asmi_sector_erase.conduit_sector_erase
			asmi_sector_protect  => asmi_sector_protect,  -- asmi_sector_protect.conduit_sector_protect
			epcq_dclk            => epcq_dclk,            --           epcq_dclk.conduit_epcq_dclk
			epcq_scein           => epcq_scein,           --          epcq_scein.conduit_epcq_scein
			epcq_sdoin           => epcq_sdoin,           --          epcq_sdoin.conduit_epcq_sdoin
			epcq_dataoe          => epcq_dataoe,          --         epcq_dataoe.conduit_epcq_dataoe
			asmi_clkin           => asmi_clkin,           --          asmi_clkin.conduit_clkin
			asmi_reset           => asmi_reset,           --          asmi_reset.conduit_reset
			asmi_sce             => asmi_sce,             --            asmi_sce.conduit_asmi_sce
			asmi_addr            => asmi_addr,            --           asmi_addr.conduit_addr
			asmi_datain          => asmi_datain,          --         asmi_datain.conduit_datain
			asmi_fast_read       => asmi_fast_read,       --      asmi_fast_read.conduit_fast_read
			asmi_rden            => asmi_rden,            --           asmi_rden.conduit_rden
			asmi_shift_bytes     => asmi_shift_bytes,     --    asmi_shift_bytes.conduit_shift_bytes
			asmi_wren            => asmi_wren,            --           asmi_wren.conduit_wren
			asmi_write           => asmi_write,           --          asmi_write.conduit_write
			asmi_rdid_out        => asmi_rdid_out,        --       asmi_rdid_out.conduit_rdid_out
			asmi_en4b_addr       => asmi_en4b_addr,       --      asmi_en4b_addr.conduit_en4b_addr
			irq                  => irq                   --    interrupt_sender.irq
		);

end architecture rtl; -- of altera_epcq_controller_core
